library verilog;
use verilog.vl_types.all;
entity simple_480p_vlg_vec_tst is
end simple_480p_vlg_vec_tst;
